program Execute_test(
    
);
    
endprogram