interface alu_if;
    logic [3:0] a_if;
    logic [3:0] b_if;
    logic [2:0] opcode_if;
    logic [3:0] result_if;
    logic carry_out_if;
    logic zero_if;
endinterface //alu_if